`default_nettype none

/////////////////////////////////////////////////////////////////
// HEADER 
//
// Module : sdreader
// Description : module to read the sd card 
// 
//
/////////////////////////////////////////////////////////////////

module sdreader (
 
);
endmodule