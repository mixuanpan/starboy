`default_nettype none

module ai_activation_unit #(
    parameter int DATA_WIDTH = 16 // bit width of feature map elements 
)(
    input logic clk, rst 
);

endmodule 