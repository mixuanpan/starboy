`timescale 1ms/10ps
module movedown_tb; 
    logic clk, rst; 
    logic [21:0][9:0][2:0] in_arr, out_arr; 
    logic [2:0] state; 
    logic [9:0] display_frame;  
    movedown mdown (.clk(clk), .rst(rst), .input_array(in_arr), .output_array(out_arr), .current_state(state)); 

    initial clk = 0; 
    always clk = #1 ~clk; 

    task tog_rst(); 
        rst = 1; #1; 
        rst = 0; 
    endtask 

    initial begin 
        $dumpfile("waves/movedown.vcd"); 
        $dumpvars(0, movedown_tb); 

        in_arr = 0; 

        // change state 
        for (integer i = 0; i <= 'd6; i++) begin 
            state = i[2:0]; 
            tog_rst();
            #5; 

            if (state == 0 || state == 'd1 || state == 'd2 || state == 'd4) begin 
                $display("output array, state: \%b", state); 
                $write("row%0d: ", 0); 
                    display_frame[0] = out_arr[0][0][1]; 
                    display_frame[1] = out_arr[0][1][1]; 
                    display_frame[2] = out_arr[0][2][1]; 
                    display_frame[3] = out_arr[0][3][1]; 
                    display_frame[4] = out_arr[0][4][1]; 
                    display_frame[5] = out_arr[0][5][1]; 
                    display_frame[6] = out_arr[0][6][1]; 
                    display_frame[7] = out_arr[0][7][1]; 
                    display_frame[8] = out_arr[0][8][1]; 
                    display_frame[9] = out_arr[0][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 1); 
                    display_frame[0] = out_arr[1][0][1]; 
                    display_frame[1] = out_arr[1][1][1]; 
                    display_frame[2] = out_arr[1][2][1]; 
                    display_frame[3] = out_arr[1][3][1]; 
                    display_frame[4] = out_arr[1][4][1]; 
                    display_frame[5] = out_arr[1][5][1]; 
                    display_frame[6] = out_arr[1][6][1]; 
                    display_frame[7] = out_arr[1][7][1]; 
                    display_frame[8] = out_arr[1][8][1]; 
                    display_frame[9] = out_arr[1][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 2); 
                    display_frame[0] = out_arr[2][0][1]; 
                    display_frame[1] = out_arr[2][1][1]; 
                    display_frame[2] = out_arr[2][2][1]; 
                    display_frame[3] = out_arr[2][3][1]; 
                    display_frame[4] = out_arr[2][4][1]; 
                    display_frame[5] = out_arr[2][5][1]; 
                    display_frame[6] = out_arr[2][6][1]; 
                    display_frame[7] = out_arr[2][7][1]; 
                    display_frame[8] = out_arr[2][8][1]; 
                    display_frame[9] = out_arr[2][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 3); 
                    display_frame[0] = out_arr[3][0][1]; 
                    display_frame[1] = out_arr[3][1][1]; 
                    display_frame[2] = out_arr[3][2][1]; 
                    display_frame[3] = out_arr[3][3][1]; 
                    display_frame[4] = out_arr[3][4][1]; 
                    display_frame[5] = out_arr[3][5][1]; 
                    display_frame[6] = out_arr[3][6][1]; 
                    display_frame[7] = out_arr[3][7][1]; 
                    display_frame[8] = out_arr[3][8][1]; 
                    display_frame[9] = out_arr[3][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 4); 
                    display_frame[0] = out_arr[4][0][1]; 
                    display_frame[1] = out_arr[4][1][1]; 
                    display_frame[2] = out_arr[4][2][1]; 
                    display_frame[3] = out_arr[4][3][1]; 
                    display_frame[4] = out_arr[4][4][1]; 
                    display_frame[5] = out_arr[4][5][1]; 
                    display_frame[6] = out_arr[4][6][1]; 
                    display_frame[7] = out_arr[4][7][1]; 
                    display_frame[8] = out_arr[4][8][1]; 
                    display_frame[9] = out_arr[4][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 5); 
                    display_frame[0] = out_arr[5][0][1]; 
                    display_frame[1] = out_arr[5][1][1]; 
                    display_frame[2] = out_arr[5][2][1]; 
                    display_frame[3] = out_arr[5][3][1]; 
                    display_frame[4] = out_arr[5][4][1]; 
                    display_frame[5] = out_arr[5][5][1]; 
                    display_frame[6] = out_arr[5][6][1]; 
                    display_frame[7] = out_arr[5][7][1]; 
                    display_frame[8] = out_arr[5][8][1]; 
                    display_frame[9] = out_arr[5][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 6); 
                    display_frame[0] = out_arr[6][0][1]; 
                    display_frame[1] = out_arr[6][1][1]; 
                    display_frame[2] = out_arr[6][2][1]; 
                    display_frame[3] = out_arr[6][3][1]; 
                    display_frame[4] = out_arr[6][4][1]; 
                    display_frame[5] = out_arr[6][5][1]; 
                    display_frame[6] = out_arr[6][6][1]; 
                    display_frame[7] = out_arr[6][7][1]; 
                    display_frame[8] = out_arr[6][8][1]; 
                    display_frame[9] = out_arr[6][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 7); 
                    display_frame[0] = out_arr[7][0][1]; 
                    display_frame[1] = out_arr[7][1][1]; 
                    display_frame[2] = out_arr[7][2][1]; 
                    display_frame[3] = out_arr[7][3][1]; 
                    display_frame[4] = out_arr[7][4][1]; 
                    display_frame[5] = out_arr[7][5][1]; 
                    display_frame[6] = out_arr[7][6][1]; 
                    display_frame[7] = out_arr[7][7][1]; 
                    display_frame[8] = out_arr[7][8][1]; 
                    display_frame[9] = out_arr[7][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 8); 
                    display_frame[0] = out_arr[8][0][1]; 
                    display_frame[1] = out_arr[8][1][1]; 
                    display_frame[2] = out_arr[8][2][1]; 
                    display_frame[3] = out_arr[8][3][1]; 
                    display_frame[4] = out_arr[8][4][1]; 
                    display_frame[5] = out_arr[8][5][1]; 
                    display_frame[6] = out_arr[8][6][1]; 
                    display_frame[7] = out_arr[8][7][1]; 
                    display_frame[8] = out_arr[8][8][1]; 
                    display_frame[9] = out_arr[8][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 9); 
                    display_frame[0] = out_arr[9][0][1]; 
                    display_frame[1] = out_arr[9][1][1]; 
                    display_frame[2] = out_arr[9][2][1]; 
                    display_frame[3] = out_arr[9][3][1]; 
                    display_frame[4] = out_arr[9][4][1]; 
                    display_frame[5] = out_arr[9][5][1]; 
                    display_frame[6] = out_arr[9][6][1]; 
                    display_frame[7] = out_arr[9][7][1]; 
                    display_frame[8] = out_arr[9][8][1]; 
                    display_frame[9] = out_arr[9][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 10); 
                    display_frame[0] = out_arr[10][0][1]; 
                    display_frame[1] = out_arr[10][1][1]; 
                    display_frame[2] = out_arr[10][2][1]; 
                    display_frame[3] = out_arr[10][3][1]; 
                    display_frame[4] = out_arr[10][4][1]; 
                    display_frame[5] = out_arr[10][5][1]; 
                    display_frame[6] = out_arr[10][6][1]; 
                    display_frame[7] = out_arr[10][7][1]; 
                    display_frame[8] = out_arr[10][8][1]; 
                    display_frame[9] = out_arr[10][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 11); 
                    display_frame[0] = out_arr[11][0][1]; 
                    display_frame[1] = out_arr[11][1][1]; 
                    display_frame[2] = out_arr[11][2][1]; 
                    display_frame[3] = out_arr[11][3][1]; 
                    display_frame[4] = out_arr[11][4][1]; 
                    display_frame[5] = out_arr[11][5][1]; 
                    display_frame[6] = out_arr[11][6][1]; 
                    display_frame[7] = out_arr[11][7][1]; 
                    display_frame[8] = out_arr[11][8][1]; 
                    display_frame[9] = out_arr[11][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 12); 
                    display_frame[0] = out_arr[12][0][1]; 
                    display_frame[1] = out_arr[12][1][1]; 
                    display_frame[2] = out_arr[12][2][1]; 
                    display_frame[3] = out_arr[12][3][1]; 
                    display_frame[4] = out_arr[12][4][1]; 
                    display_frame[5] = out_arr[12][5][1]; 
                    display_frame[6] = out_arr[12][6][1]; 
                    display_frame[7] = out_arr[12][7][1]; 
                    display_frame[8] = out_arr[12][8][1]; 
                    display_frame[9] = out_arr[12][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 13); 
                    display_frame[0] = out_arr[13][0][1]; 
                    display_frame[1] = out_arr[13][1][1]; 
                    display_frame[2] = out_arr[13][2][1]; 
                    display_frame[3] = out_arr[13][3][1]; 
                    display_frame[4] = out_arr[13][4][1]; 
                    display_frame[5] = out_arr[13][5][1]; 
                    display_frame[6] = out_arr[13][6][1]; 
                    display_frame[7] = out_arr[13][7][1]; 
                    display_frame[8] = out_arr[13][8][1]; 
                    display_frame[9] = out_arr[13][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 14); 
                    display_frame[0] = out_arr[14][0][1]; 
                    display_frame[1] = out_arr[14][1][1]; 
                    display_frame[2] = out_arr[14][2][1]; 
                    display_frame[3] = out_arr[14][3][1]; 
                    display_frame[4] = out_arr[14][4][1]; 
                    display_frame[5] = out_arr[14][5][1]; 
                    display_frame[6] = out_arr[14][6][1]; 
                    display_frame[7] = out_arr[14][7][1]; 
                    display_frame[8] = out_arr[14][8][1]; 
                    display_frame[9] = out_arr[14][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 15); 
                    display_frame[0] = out_arr[15][0][1]; 
                    display_frame[1] = out_arr[15][1][1]; 
                    display_frame[2] = out_arr[15][2][1]; 
                    display_frame[3] = out_arr[15][3][1]; 
                    display_frame[4] = out_arr[15][4][1]; 
                    display_frame[5] = out_arr[15][5][1]; 
                    display_frame[6] = out_arr[15][6][1]; 
                    display_frame[7] = out_arr[15][7][1]; 
                    display_frame[8] = out_arr[15][8][1]; 
                    display_frame[9] = out_arr[15][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 16); 
                    display_frame[0] = out_arr[16][0][1]; 
                    display_frame[1] = out_arr[16][1][1]; 
                    display_frame[2] = out_arr[16][2][1]; 
                    display_frame[3] = out_arr[16][3][1]; 
                    display_frame[4] = out_arr[16][4][1]; 
                    display_frame[5] = out_arr[16][5][1]; 
                    display_frame[6] = out_arr[16][6][1]; 
                    display_frame[7] = out_arr[16][7][1]; 
                    display_frame[8] = out_arr[16][8][1]; 
                    display_frame[9] = out_arr[16][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 17); 
                    display_frame[0] = out_arr[17][0][1]; 
                    display_frame[1] = out_arr[17][1][1]; 
                    display_frame[2] = out_arr[17][2][1]; 
                    display_frame[3] = out_arr[17][3][1]; 
                    display_frame[4] = out_arr[17][4][1]; 
                    display_frame[5] = out_arr[17][5][1]; 
                    display_frame[6] = out_arr[17][6][1]; 
                    display_frame[7] = out_arr[17][7][1]; 
                    display_frame[8] = out_arr[17][8][1]; 
                    display_frame[9] = out_arr[17][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 18); 
                    display_frame[0] = out_arr[18][0][1]; 
                    display_frame[1] = out_arr[18][1][1]; 
                    display_frame[2] = out_arr[18][2][1]; 
                    display_frame[3] = out_arr[18][3][1]; 
                    display_frame[4] = out_arr[18][4][1]; 
                    display_frame[5] = out_arr[18][5][1]; 
                    display_frame[6] = out_arr[18][6][1]; 
                    display_frame[7] = out_arr[18][7][1]; 
                    display_frame[8] = out_arr[18][8][1]; 
                    display_frame[9] = out_arr[18][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 19); 
                    display_frame[0] = out_arr[19][0][1]; 
                    display_frame[1] = out_arr[19][1][1]; 
                    display_frame[2] = out_arr[19][2][1]; 
                    display_frame[3] = out_arr[19][3][1]; 
                    display_frame[4] = out_arr[19][4][1]; 
                    display_frame[5] = out_arr[19][5][1]; 
                    display_frame[6] = out_arr[19][6][1]; 
                    display_frame[7] = out_arr[19][7][1]; 
                    display_frame[8] = out_arr[19][8][1]; 
                    display_frame[9] = out_arr[19][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 20); 
                    display_frame[0] = out_arr[20][0][1]; 
                    display_frame[1] = out_arr[20][1][1]; 
                    display_frame[2] = out_arr[20][2][1]; 
                    display_frame[3] = out_arr[20][3][1]; 
                    display_frame[4] = out_arr[20][4][1]; 
                    display_frame[5] = out_arr[20][5][1]; 
                    display_frame[6] = out_arr[20][6][1]; 
                    display_frame[7] = out_arr[20][7][1]; 
                    display_frame[8] = out_arr[20][8][1]; 
                    display_frame[9] = out_arr[20][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 21); 
                    display_frame[0] = out_arr[21][0][1]; 
                    display_frame[1] = out_arr[21][1][1]; 
                    display_frame[2] = out_arr[21][2][1]; 
                    display_frame[3] = out_arr[21][3][1]; 
                    display_frame[4] = out_arr[21][4][1]; 
                    display_frame[5] = out_arr[21][5][1]; 
                    display_frame[6] = out_arr[21][6][1]; 
                    display_frame[7] = out_arr[21][7][1]; 
                    display_frame[8] = out_arr[21][8][1]; 
                    display_frame[9] = out_arr[21][9][1]; 
                $write("%b", display_frame); 
                $write("\n"); 
            end else if (state == 'd3) begin 
                $write("row%0d: ", 0); 
                    display_frame[0] = out_arr[0][0][0]; 
                    display_frame[1] = out_arr[0][1][0]; 
                    display_frame[2] = out_arr[0][2][0]; 
                    display_frame[3] = out_arr[0][3][0]; 
                    display_frame[4] = out_arr[0][4][0]; 
                    display_frame[5] = out_arr[0][5][0]; 
                    display_frame[6] = out_arr[0][6][0]; 
                    display_frame[7] = out_arr[0][7][0]; 
                    display_frame[8] = out_arr[0][8][0]; 
                    display_frame[9] = out_arr[0][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 1); 
                    display_frame[0] = out_arr[1][0][0]; 
                    display_frame[1] = out_arr[1][1][0]; 
                    display_frame[2] = out_arr[1][2][0]; 
                    display_frame[3] = out_arr[1][3][0]; 
                    display_frame[4] = out_arr[1][4][0]; 
                    display_frame[5] = out_arr[1][5][0]; 
                    display_frame[6] = out_arr[1][6][0]; 
                    display_frame[7] = out_arr[1][7][0]; 
                    display_frame[8] = out_arr[1][8][0]; 
                    display_frame[9] = out_arr[1][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 2); 
                    display_frame[0] = out_arr[2][0][0]; 
                    display_frame[1] = out_arr[2][1][0]; 
                    display_frame[2] = out_arr[2][2][0]; 
                    display_frame[3] = out_arr[2][3][0]; 
                    display_frame[4] = out_arr[2][4][0]; 
                    display_frame[5] = out_arr[2][5][0]; 
                    display_frame[6] = out_arr[2][6][0]; 
                    display_frame[7] = out_arr[2][7][0]; 
                    display_frame[8] = out_arr[2][8][0]; 
                    display_frame[9] = out_arr[2][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 3); 
                    display_frame[0] = out_arr[3][0][0]; 
                    display_frame[1] = out_arr[3][1][0]; 
                    display_frame[2] = out_arr[3][2][0]; 
                    display_frame[3] = out_arr[3][3][0]; 
                    display_frame[4] = out_arr[3][4][0]; 
                    display_frame[5] = out_arr[3][5][0]; 
                    display_frame[6] = out_arr[3][6][0]; 
                    display_frame[7] = out_arr[3][7][0]; 
                    display_frame[8] = out_arr[3][8][0]; 
                    display_frame[9] = out_arr[3][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 4); 
                    display_frame[0] = out_arr[4][0][0]; 
                    display_frame[1] = out_arr[4][1][0]; 
                    display_frame[2] = out_arr[4][2][0]; 
                    display_frame[3] = out_arr[4][3][0]; 
                    display_frame[4] = out_arr[4][4][0]; 
                    display_frame[5] = out_arr[4][5][0]; 
                    display_frame[6] = out_arr[4][6][0]; 
                    display_frame[7] = out_arr[4][7][0]; 
                    display_frame[8] = out_arr[4][8][0]; 
                    display_frame[9] = out_arr[4][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 5); 
                    display_frame[0] = out_arr[5][0][0]; 
                    display_frame[1] = out_arr[5][1][0]; 
                    display_frame[2] = out_arr[5][2][0]; 
                    display_frame[3] = out_arr[5][3][0]; 
                    display_frame[4] = out_arr[5][4][0]; 
                    display_frame[5] = out_arr[5][5][0]; 
                    display_frame[6] = out_arr[5][6][0]; 
                    display_frame[7] = out_arr[5][7][0]; 
                    display_frame[8] = out_arr[5][8][0]; 
                    display_frame[9] = out_arr[5][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 6); 
                    display_frame[0] = out_arr[6][0][0]; 
                    display_frame[1] = out_arr[6][1][0]; 
                    display_frame[2] = out_arr[6][2][0]; 
                    display_frame[3] = out_arr[6][3][0]; 
                    display_frame[4] = out_arr[6][4][0]; 
                    display_frame[5] = out_arr[6][5][0]; 
                    display_frame[6] = out_arr[6][6][0]; 
                    display_frame[7] = out_arr[6][7][0]; 
                    display_frame[8] = out_arr[6][8][0]; 
                    display_frame[9] = out_arr[6][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 7); 
                    display_frame[0] = out_arr[7][0][0]; 
                    display_frame[1] = out_arr[7][1][0]; 
                    display_frame[2] = out_arr[7][2][0]; 
                    display_frame[3] = out_arr[7][3][0]; 
                    display_frame[4] = out_arr[7][4][0]; 
                    display_frame[5] = out_arr[7][5][0]; 
                    display_frame[6] = out_arr[7][6][0]; 
                    display_frame[7] = out_arr[7][7][0]; 
                    display_frame[8] = out_arr[7][8][0]; 
                    display_frame[9] = out_arr[7][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 8); 
                    display_frame[0] = out_arr[8][0][0]; 
                    display_frame[1] = out_arr[8][1][0]; 
                    display_frame[2] = out_arr[8][2][0]; 
                    display_frame[3] = out_arr[8][3][0]; 
                    display_frame[4] = out_arr[8][4][0]; 
                    display_frame[5] = out_arr[8][5][0]; 
                    display_frame[6] = out_arr[8][6][0]; 
                    display_frame[7] = out_arr[8][7][0]; 
                    display_frame[8] = out_arr[8][8][0]; 
                    display_frame[9] = out_arr[8][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 9); 
                    display_frame[0] = out_arr[9][0][0]; 
                    display_frame[1] = out_arr[9][1][0]; 
                    display_frame[2] = out_arr[9][2][0]; 
                    display_frame[3] = out_arr[9][3][0]; 
                    display_frame[4] = out_arr[9][4][0]; 
                    display_frame[5] = out_arr[9][5][0]; 
                    display_frame[6] = out_arr[9][6][0]; 
                    display_frame[7] = out_arr[9][7][0]; 
                    display_frame[8] = out_arr[9][8][0]; 
                    display_frame[9] = out_arr[9][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 10); 
                    display_frame[0] = out_arr[10][0][0]; 
                    display_frame[1] = out_arr[10][1][0]; 
                    display_frame[2] = out_arr[10][2][0]; 
                    display_frame[3] = out_arr[10][3][0]; 
                    display_frame[4] = out_arr[10][4][0]; 
                    display_frame[5] = out_arr[10][5][0]; 
                    display_frame[6] = out_arr[10][6][0]; 
                    display_frame[7] = out_arr[10][7][0]; 
                    display_frame[8] = out_arr[10][8][0]; 
                    display_frame[9] = out_arr[10][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 11); 
                    display_frame[0] = out_arr[11][0][0]; 
                    display_frame[1] = out_arr[11][1][0]; 
                    display_frame[2] = out_arr[11][2][0]; 
                    display_frame[3] = out_arr[11][3][0]; 
                    display_frame[4] = out_arr[11][4][0]; 
                    display_frame[5] = out_arr[11][5][0]; 
                    display_frame[6] = out_arr[11][6][0]; 
                    display_frame[7] = out_arr[11][7][0]; 
                    display_frame[8] = out_arr[11][8][0]; 
                    display_frame[9] = out_arr[11][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 12); 
                    display_frame[0] = out_arr[12][0][0]; 
                    display_frame[1] = out_arr[12][1][0]; 
                    display_frame[2] = out_arr[12][2][0]; 
                    display_frame[3] = out_arr[12][3][0]; 
                    display_frame[4] = out_arr[12][4][0]; 
                    display_frame[5] = out_arr[12][5][0]; 
                    display_frame[6] = out_arr[12][6][0]; 
                    display_frame[7] = out_arr[12][7][0]; 
                    display_frame[8] = out_arr[12][8][0]; 
                    display_frame[9] = out_arr[12][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 13); 
                    display_frame[0] = out_arr[13][0][0]; 
                    display_frame[1] = out_arr[13][1][0]; 
                    display_frame[2] = out_arr[13][2][0]; 
                    display_frame[3] = out_arr[13][3][0]; 
                    display_frame[4] = out_arr[13][4][0]; 
                    display_frame[5] = out_arr[13][5][0]; 
                    display_frame[6] = out_arr[13][6][0]; 
                    display_frame[7] = out_arr[13][7][0]; 
                    display_frame[8] = out_arr[13][8][0]; 
                    display_frame[9] = out_arr[13][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 14); 
                    display_frame[0] = out_arr[14][0][0]; 
                    display_frame[1] = out_arr[14][1][0]; 
                    display_frame[2] = out_arr[14][2][0]; 
                    display_frame[3] = out_arr[14][3][0]; 
                    display_frame[4] = out_arr[14][4][0]; 
                    display_frame[5] = out_arr[14][5][0]; 
                    display_frame[6] = out_arr[14][6][0]; 
                    display_frame[7] = out_arr[14][7][0]; 
                    display_frame[8] = out_arr[14][8][0]; 
                    display_frame[9] = out_arr[14][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 15); 
                    display_frame[0] = out_arr[15][0][0]; 
                    display_frame[1] = out_arr[15][1][0]; 
                    display_frame[2] = out_arr[15][2][0]; 
                    display_frame[3] = out_arr[15][3][0]; 
                    display_frame[4] = out_arr[15][4][0]; 
                    display_frame[5] = out_arr[15][5][0]; 
                    display_frame[6] = out_arr[15][6][0]; 
                    display_frame[7] = out_arr[15][7][0]; 
                    display_frame[8] = out_arr[15][8][0]; 
                    display_frame[9] = out_arr[15][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 16); 
                    display_frame[0] = out_arr[16][0][0]; 
                    display_frame[1] = out_arr[16][1][0]; 
                    display_frame[2] = out_arr[16][2][0]; 
                    display_frame[3] = out_arr[16][3][0]; 
                    display_frame[4] = out_arr[16][4][0]; 
                    display_frame[5] = out_arr[16][5][0]; 
                    display_frame[6] = out_arr[16][6][0]; 
                    display_frame[7] = out_arr[16][7][0]; 
                    display_frame[8] = out_arr[16][8][0]; 
                    display_frame[9] = out_arr[16][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 17); 
                    display_frame[0] = out_arr[17][0][0]; 
                    display_frame[1] = out_arr[17][1][0]; 
                    display_frame[2] = out_arr[17][2][0]; 
                    display_frame[3] = out_arr[17][3][0]; 
                    display_frame[4] = out_arr[17][4][0]; 
                    display_frame[5] = out_arr[17][5][0]; 
                    display_frame[6] = out_arr[17][6][0]; 
                    display_frame[7] = out_arr[17][7][0]; 
                    display_frame[8] = out_arr[17][8][0]; 
                    display_frame[9] = out_arr[17][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 18); 
                    display_frame[0] = out_arr[18][0][0]; 
                    display_frame[1] = out_arr[18][1][0]; 
                    display_frame[2] = out_arr[18][2][0]; 
                    display_frame[3] = out_arr[18][3][0]; 
                    display_frame[4] = out_arr[18][4][0]; 
                    display_frame[5] = out_arr[18][5][0]; 
                    display_frame[6] = out_arr[18][6][0]; 
                    display_frame[7] = out_arr[18][7][0]; 
                    display_frame[8] = out_arr[18][8][0]; 
                    display_frame[9] = out_arr[18][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 19); 
                    display_frame[0] = out_arr[19][0][0]; 
                    display_frame[1] = out_arr[19][1][0]; 
                    display_frame[2] = out_arr[19][2][0]; 
                    display_frame[3] = out_arr[19][3][0]; 
                    display_frame[4] = out_arr[19][4][0]; 
                    display_frame[5] = out_arr[19][5][0]; 
                    display_frame[6] = out_arr[19][6][0]; 
                    display_frame[7] = out_arr[19][7][0]; 
                    display_frame[8] = out_arr[19][8][0]; 
                    display_frame[9] = out_arr[19][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 20); 
                    display_frame[0] = out_arr[20][0][0]; 
                    display_frame[1] = out_arr[20][1][0]; 
                    display_frame[2] = out_arr[20][2][0]; 
                    display_frame[3] = out_arr[20][3][0]; 
                    display_frame[4] = out_arr[20][4][0]; 
                    display_frame[5] = out_arr[20][5][0]; 
                    display_frame[6] = out_arr[20][6][0]; 
                    display_frame[7] = out_arr[20][7][0]; 
                    display_frame[8] = out_arr[20][8][0]; 
                    display_frame[9] = out_arr[20][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 

                $write("row%0d: ", 21); 
                    display_frame[0] = out_arr[21][0][0]; 
                    display_frame[1] = out_arr[21][1][0]; 
                    display_frame[2] = out_arr[21][2][0]; 
                    display_frame[3] = out_arr[21][3][0]; 
                    display_frame[4] = out_arr[21][4][0]; 
                    display_frame[5] = out_arr[21][5][0]; 
                    display_frame[6] = out_arr[21][6][0]; 
                    display_frame[7] = out_arr[21][7][0]; 
                    display_frame[8] = out_arr[21][8][0]; 
                    display_frame[9] = out_arr[21][9][0]; 
                $write("%b", display_frame); 
                $write("\n"); 
            end else begin 
                $write("row%0d: ", 0); 
                display_frame[0] = out_arr[0][0][2]; 
                display_frame[1] = out_arr[0][1][2]; 
                display_frame[2] = out_arr[0][2][2]; 
                display_frame[3] = out_arr[0][3][2]; 
                display_frame[4] = out_arr[0][4][2]; 
                display_frame[5] = out_arr[0][5][2]; 
                display_frame[6] = out_arr[0][6][2]; 
                display_frame[7] = out_arr[0][7][2]; 
                display_frame[8] = out_arr[0][8][2]; 
                display_frame[9] = out_arr[0][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 1); 
                display_frame[0] = out_arr[1][0][2]; 
                display_frame[1] = out_arr[1][1][2]; 
                display_frame[2] = out_arr[1][2][2]; 
                display_frame[3] = out_arr[1][3][2]; 
                display_frame[4] = out_arr[1][4][2]; 
                display_frame[5] = out_arr[1][5][2]; 
                display_frame[6] = out_arr[1][6][2]; 
                display_frame[7] = out_arr[1][7][2]; 
                display_frame[8] = out_arr[1][8][2]; 
                display_frame[9] = out_arr[1][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 2); 
                display_frame[0] = out_arr[2][0][2]; 
                display_frame[1] = out_arr[2][1][2]; 
                display_frame[2] = out_arr[2][2][2]; 
                display_frame[3] = out_arr[2][3][2]; 
                display_frame[4] = out_arr[2][4][2]; 
                display_frame[5] = out_arr[2][5][2]; 
                display_frame[6] = out_arr[2][6][2]; 
                display_frame[7] = out_arr[2][7][2]; 
                display_frame[8] = out_arr[2][8][2]; 
                display_frame[9] = out_arr[2][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 3); 
                display_frame[0] = out_arr[3][0][2]; 
                display_frame[1] = out_arr[3][1][2]; 
                display_frame[2] = out_arr[3][2][2]; 
                display_frame[3] = out_arr[3][3][2]; 
                display_frame[4] = out_arr[3][4][2]; 
                display_frame[5] = out_arr[3][5][2]; 
                display_frame[6] = out_arr[3][6][2]; 
                display_frame[7] = out_arr[3][7][2]; 
                display_frame[8] = out_arr[3][8][2]; 
                display_frame[9] = out_arr[3][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 4); 
                display_frame[0] = out_arr[4][0][2]; 
                display_frame[1] = out_arr[4][1][2]; 
                display_frame[2] = out_arr[4][2][2]; 
                display_frame[3] = out_arr[4][3][2]; 
                display_frame[4] = out_arr[4][4][2]; 
                display_frame[5] = out_arr[4][5][2]; 
                display_frame[6] = out_arr[4][6][2]; 
                display_frame[7] = out_arr[4][7][2]; 
                display_frame[8] = out_arr[4][8][2]; 
                display_frame[9] = out_arr[4][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 5); 
                display_frame[0] = out_arr[5][0][2]; 
                display_frame[1] = out_arr[5][1][2]; 
                display_frame[2] = out_arr[5][2][2]; 
                display_frame[3] = out_arr[5][3][2]; 
                display_frame[4] = out_arr[5][4][2]; 
                display_frame[5] = out_arr[5][5][2]; 
                display_frame[6] = out_arr[5][6][2]; 
                display_frame[7] = out_arr[5][7][2]; 
                display_frame[8] = out_arr[5][8][2]; 
                display_frame[9] = out_arr[5][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 6); 
                display_frame[0] = out_arr[6][0][2]; 
                display_frame[1] = out_arr[6][1][2]; 
                display_frame[2] = out_arr[6][2][2]; 
                display_frame[3] = out_arr[6][3][2]; 
                display_frame[4] = out_arr[6][4][2]; 
                display_frame[5] = out_arr[6][5][2]; 
                display_frame[6] = out_arr[6][6][2]; 
                display_frame[7] = out_arr[6][7][2]; 
                display_frame[8] = out_arr[6][8][2]; 
                display_frame[9] = out_arr[6][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 7); 
                display_frame[0] = out_arr[7][0][2]; 
                display_frame[1] = out_arr[7][1][2]; 
                display_frame[2] = out_arr[7][2][2]; 
                display_frame[3] = out_arr[7][3][2]; 
                display_frame[4] = out_arr[7][4][2]; 
                display_frame[5] = out_arr[7][5][2]; 
                display_frame[6] = out_arr[7][6][2]; 
                display_frame[7] = out_arr[7][7][2]; 
                display_frame[8] = out_arr[7][8][2]; 
                display_frame[9] = out_arr[7][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 8); 
                display_frame[0] = out_arr[8][0][2]; 
                display_frame[1] = out_arr[8][1][2]; 
                display_frame[2] = out_arr[8][2][2]; 
                display_frame[3] = out_arr[8][3][2]; 
                display_frame[4] = out_arr[8][4][2]; 
                display_frame[5] = out_arr[8][5][2]; 
                display_frame[6] = out_arr[8][6][2]; 
                display_frame[7] = out_arr[8][7][2]; 
                display_frame[8] = out_arr[8][8][2]; 
                display_frame[9] = out_arr[8][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 9); 
                display_frame[0] = out_arr[9][0][2]; 
                display_frame[1] = out_arr[9][1][2]; 
                display_frame[2] = out_arr[9][2][2]; 
                display_frame[3] = out_arr[9][3][2]; 
                display_frame[4] = out_arr[9][4][2]; 
                display_frame[5] = out_arr[9][5][2]; 
                display_frame[6] = out_arr[9][6][2]; 
                display_frame[7] = out_arr[9][7][2]; 
                display_frame[8] = out_arr[9][8][2]; 
                display_frame[9] = out_arr[9][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 10); 
                display_frame[0] = out_arr[10][0][2]; 
                display_frame[1] = out_arr[10][1][2]; 
                display_frame[2] = out_arr[10][2][2]; 
                display_frame[3] = out_arr[10][3][2]; 
                display_frame[4] = out_arr[10][4][2]; 
                display_frame[5] = out_arr[10][5][2]; 
                display_frame[6] = out_arr[10][6][2]; 
                display_frame[7] = out_arr[10][7][2]; 
                display_frame[8] = out_arr[10][8][2]; 
                display_frame[9] = out_arr[10][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 11); 
                display_frame[0] = out_arr[11][0][2]; 
                display_frame[1] = out_arr[11][1][2]; 
                display_frame[2] = out_arr[11][2][2]; 
                display_frame[3] = out_arr[11][3][2]; 
                display_frame[4] = out_arr[11][4][2]; 
                display_frame[5] = out_arr[11][5][2]; 
                display_frame[6] = out_arr[11][6][2]; 
                display_frame[7] = out_arr[11][7][2]; 
                display_frame[8] = out_arr[11][8][2]; 
                display_frame[9] = out_arr[11][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 12); 
                display_frame[0] = out_arr[12][0][2]; 
                display_frame[1] = out_arr[12][1][2]; 
                display_frame[2] = out_arr[12][2][2]; 
                display_frame[3] = out_arr[12][3][2]; 
                display_frame[4] = out_arr[12][4][2]; 
                display_frame[5] = out_arr[12][5][2]; 
                display_frame[6] = out_arr[12][6][2]; 
                display_frame[7] = out_arr[12][7][2]; 
                display_frame[8] = out_arr[12][8][2]; 
                display_frame[9] = out_arr[12][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 13); 
                display_frame[0] = out_arr[13][0][2]; 
                display_frame[1] = out_arr[13][1][2]; 
                display_frame[2] = out_arr[13][2][2]; 
                display_frame[3] = out_arr[13][3][2]; 
                display_frame[4] = out_arr[13][4][2]; 
                display_frame[5] = out_arr[13][5][2]; 
                display_frame[6] = out_arr[13][6][2]; 
                display_frame[7] = out_arr[13][7][2]; 
                display_frame[8] = out_arr[13][8][2]; 
                display_frame[9] = out_arr[13][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 14); 
                display_frame[0] = out_arr[14][0][2]; 
                display_frame[1] = out_arr[14][1][2]; 
                display_frame[2] = out_arr[14][2][2]; 
                display_frame[3] = out_arr[14][3][2]; 
                display_frame[4] = out_arr[14][4][2]; 
                display_frame[5] = out_arr[14][5][2]; 
                display_frame[6] = out_arr[14][6][2]; 
                display_frame[7] = out_arr[14][7][2]; 
                display_frame[8] = out_arr[14][8][2]; 
                display_frame[9] = out_arr[14][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 15); 
                display_frame[0] = out_arr[15][0][2]; 
                display_frame[1] = out_arr[15][1][2]; 
                display_frame[2] = out_arr[15][2][2]; 
                display_frame[3] = out_arr[15][3][2]; 
                display_frame[4] = out_arr[15][4][2]; 
                display_frame[5] = out_arr[15][5][2]; 
                display_frame[6] = out_arr[15][6][2]; 
                display_frame[7] = out_arr[15][7][2]; 
                display_frame[8] = out_arr[15][8][2]; 
                display_frame[9] = out_arr[15][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 16); 
                display_frame[0] = out_arr[16][0][2]; 
                display_frame[1] = out_arr[16][1][2]; 
                display_frame[2] = out_arr[16][2][2]; 
                display_frame[3] = out_arr[16][3][2]; 
                display_frame[4] = out_arr[16][4][2]; 
                display_frame[5] = out_arr[16][5][2]; 
                display_frame[6] = out_arr[16][6][2]; 
                display_frame[7] = out_arr[16][7][2]; 
                display_frame[8] = out_arr[16][8][2]; 
                display_frame[9] = out_arr[16][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 17); 
                display_frame[0] = out_arr[17][0][2]; 
                display_frame[1] = out_arr[17][1][2]; 
                display_frame[2] = out_arr[17][2][2]; 
                display_frame[3] = out_arr[17][3][2]; 
                display_frame[4] = out_arr[17][4][2]; 
                display_frame[5] = out_arr[17][5][2]; 
                display_frame[6] = out_arr[17][6][2]; 
                display_frame[7] = out_arr[17][7][2]; 
                display_frame[8] = out_arr[17][8][2]; 
                display_frame[9] = out_arr[17][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 18); 
                display_frame[0] = out_arr[18][0][2]; 
                display_frame[1] = out_arr[18][1][2]; 
                display_frame[2] = out_arr[18][2][2]; 
                display_frame[3] = out_arr[18][3][2]; 
                display_frame[4] = out_arr[18][4][2]; 
                display_frame[5] = out_arr[18][5][2]; 
                display_frame[6] = out_arr[18][6][2]; 
                display_frame[7] = out_arr[18][7][2]; 
                display_frame[8] = out_arr[18][8][2]; 
                display_frame[9] = out_arr[18][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 19); 
                display_frame[0] = out_arr[19][0][2]; 
                display_frame[1] = out_arr[19][1][2]; 
                display_frame[2] = out_arr[19][2][2]; 
                display_frame[3] = out_arr[19][3][2]; 
                display_frame[4] = out_arr[19][4][2]; 
                display_frame[5] = out_arr[19][5][2]; 
                display_frame[6] = out_arr[19][6][2]; 
                display_frame[7] = out_arr[19][7][2]; 
                display_frame[8] = out_arr[19][8][2]; 
                display_frame[9] = out_arr[19][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 20); 
                display_frame[0] = out_arr[20][0][2]; 
                display_frame[1] = out_arr[20][1][2]; 
                display_frame[2] = out_arr[20][2][2]; 
                display_frame[3] = out_arr[20][3][2]; 
                display_frame[4] = out_arr[20][4][2]; 
                display_frame[5] = out_arr[20][5][2]; 
                display_frame[6] = out_arr[20][6][2]; 
                display_frame[7] = out_arr[20][7][2]; 
                display_frame[8] = out_arr[20][8][2]; 
                display_frame[9] = out_arr[20][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            $write("row%0d: ", 21); 
                display_frame[0] = out_arr[21][0][2]; 
                display_frame[1] = out_arr[21][1][2]; 
                display_frame[2] = out_arr[21][2][2]; 
                display_frame[3] = out_arr[21][3][2]; 
                display_frame[4] = out_arr[21][4][2]; 
                display_frame[5] = out_arr[21][5][2]; 
                display_frame[6] = out_arr[21][6][2]; 
                display_frame[7] = out_arr[21][7][2]; 
                display_frame[8] = out_arr[21][8][2]; 
                display_frame[9] = out_arr[21][9][2]; 
            $write("%b", display_frame); 
            $write("\n"); 

            end
        end


    end
endmodule 