`default_nettype none
module read_block (
  //put your ports here
);
//your code starts here ...
endmodule