module frameBuffer(

);

//buff men
endmodule