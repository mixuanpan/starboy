module iloveplayer333(
    input logic myles
    input logic querimit
);



assign fix fix 
endmodule