`default_nettype none
/////////////////////////////////////////////////////////////////
// HEADER 
//
// Module : ai_mc_rd_arbiter   
// Description : Reads out the Output Feature-Map BRAM for write-back
//               Instantiates an Address Generator to step through the OFM, 
//               then pulls data from the ofm_buffer and presents it as a
//                valid-ready stream to the write-FIFO / serializer. 
//
/////////////////////////////////////////////////////////////////
module ai_mc_rd_arbiter (
    parameter int ADDR_W = 32, // bits of the ofm address 
    parameter int LEN_W = 16, // width of the length (in beats)
    parameter int  DATA_W = 32 // width of each word 
)(
    input logic clk, rst, 
    
);

endmodule 