<<<<<<< HEAD
`default_nettype none
/////////////////////////////////////////////////////////////////
// HEADER 
//
// Module : collision  
// Description : tetris collision logic  
// 
//
/////////////////////////////////////////////////////////////////
module collision (
    input logic [4:0] blockY, 
    input logic [3:0] blockX, 
    input logic [3:0][3:0] current_block_pattern, 
    input logic [19:0][9:0] stored_array, 
    output collision_bottom, collision_left, collision_right, 
    output logic [19:0][9:0] falling_block_display
);

    logic [4:0] row_ext;
    logic [3:0] col_ext;
    logic [4:0] abs_row;
    logic [3:0] abs_col;

    //collision logic
    always_comb begin
        collision_bottom       = 1'b0;
        collision_left         = 1'b0;
        collision_right        = 1'b0;
        falling_block_display  = '0;

        // 4×4 nested loop over the current tetromino pattern
        for (int row = 0; row < 4; row++) begin
            for (int col = 0; col < 4; col++) begin
                row_ext = {3'b000, row[1:0]}; 
                col_ext = {2'b00, col[1:0]}; 

                abs_row = blockY + row_ext; 
                abs_col = blockX + col_ext;

                if (current_block_pattern[row][col]) begin
                    // draw the pixel
                    if (abs_row < 5'd20 && abs_col < 4'd10) begin 
                        falling_block_display[abs_row][abs_col] = 1'b1;        
                    end 
                    // bottom collision
                    if (abs_row + 1 >= 5'd20 ||
                    ((abs_row + 1) < 5'd20 &&
                        stored_array[abs_row + 1][abs_col]))
                        collision_bottom = 1'b1;

                    // left collision
                    if (abs_col == 0 ||
                    (abs_col > 0 && stored_array[abs_row][abs_col - 1]))
                        collision_left = 1'b1;

                    // right collision
                    if (abs_col + 1 >= 4'd10 ||
                    ((abs_col + 1) < 4'd10 &&
                        stored_array[abs_row][abs_col + 1]))
                        collision_right = 1'b1;
                end
            end
        end
    end
endmodule 
=======
module collision (
    input logic [4:0] blockY,
    input logic [3:0] blockX,
    input logic [3:0][3:0] current_block_pattern,
    input logic [19:0][9:0] stored_array,
    output logic collision_bottom,
    output logic collision_left,
    output logic collision_right,
    output logic [19:0][9:0] falling_block_display
);

logic [4:0] row_ext;
logic [3:0] col_ext;
logic [4:0] abs_row;
logic [3:0] abs_col;

// Collision logic and display generation
always_comb begin
    collision_bottom = 1'b0;
    collision_left = 1'b0;
    collision_right = 1'b0;
    falling_block_display = '0;

    for (int row = 0; row < 4; row++) begin
        for (int col = 0; col < 4; col++) begin
            row_ext = {3'b000, row[1:0]}; 
            col_ext = {2'b00, col[1:0]}; 

            abs_row = blockY + row_ext; 
            abs_col = blockX + col_ext;

            if (current_block_pattern[row][col]) begin
                if (abs_row < 5'd20 && abs_col < 4'd10) begin 
                    falling_block_display[abs_row][abs_col] = 1'b1;        
                end 
                
                if (abs_row + 1 >= 5'd20 ||
                   ((abs_row + 1) < 5'd20 &&
                    stored_array[abs_row + 1][abs_col]))
                    collision_bottom = 1'b1;

                if (abs_col == 0 ||
                   (abs_col > 0 && stored_array[abs_row][abs_col - 1]))
                    collision_left = 1'b1;

                if (abs_col + 1 >= 4'd10 ||
                   ((abs_col + 1) < 4'd10 &&
                    stored_array[abs_row][abs_col + 1]))
                    collision_right = 1'b1;
            end
        end
    end
end

endmodule
>>>>>>> 021eefa44bd0c4666ebf66705ed9f98d3ea607ec
