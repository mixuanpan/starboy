// `timescale 1ms/10ps
// module ai_cu_id_tb(

// )