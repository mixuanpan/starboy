`default_nettype none
module fa (
  //put your ports here
);
//your code starts here ...
endmodule