module iloveplayer333(
    input logic myles
    input logic querimit
);

endmodule