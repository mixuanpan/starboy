`default_nettype none

/////////////////////////////////////////////////////////////////
// HEADER 
//
// Module : inputbus
// Description : converts the pb inputs to moves
// 
//
/////////////////////////////////////////////////////////////////

module inputbus (
  input logic [3:0] in, 
  input logic enable, 
  output logic [7:0] out
);

endmodule