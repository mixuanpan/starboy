//gurt
