`default_nettype none 
/////////////////////////////////////////////////////////////////
// HEADER 
//
// Module : clkdiv1hz
// Description : takes 25mhz clock and turns it into 1 hz, subject to change
// 
//
/////////////////////////////////////////////////////////////////

im workign on this rn